entity SystemE is
  port (A,B,C : in bit;
        F: out bit);
end entity;
  
architecture SystemE_arch of SystemE is
  
  signal An, Bn, Cn : bit;
  signal m1, m3, m4, m6 : bit;

  begin
    An <= not A;
    Bn <= not B;
    Cn <= not C;

    m1 <= An and Bn and C;
    m3 <= An and B and C;
    m4 <= A and Bn and Cn;
    m6 <= A and B and Cn;

    F <= m1 or m3 or m4 or m6;

end architecture;
